/**
 * Configuration Registers
 * 
 * Description:
 *   Stores configuration parameters for the PE Controller.
 *   Accessible via a simple 32-bit register interface.
 *
 * Address Map:
 *   0x00: Control Register
 *         Bit 0: Start (RW, Auto-clears or Pulse?) -> Let's make it a pulse generator or level.
 *                Controller expects a 'start' signal.
 *   0x04: Status Register (RO)
 *         Bit 0: Done
 *   0x08: Kernel Dimensions
 *         Bits 3:0   -> Kernel Width (KW)
 *         Bits 7:4   -> Reserved
 *         Bits 11:8  -> Kernel Height (KH)
 *   0x0C: Input Dimensions
 *         Bits 7:0   -> Input Width (W)
 *         Bits 15:8  -> Input Height (H)
 *   0x10: Stride & Padding
 *         Bits 3:0   -> Stride
 *         Bits 7:4   -> Padding
 *   0x14: Output Dimensions
 *         Bits 7:0   -> Output Width
 *         Bits 15:8  -> Output Height
 *   0x18: Channel Configuration
 *         Bits 7:0   -> Input Channels (must be 16 or multiple of 16)
 *         Bits 15:8  -> Output Channels (Total, auto-batched in groups of 16)
 *
 * Author: shealligh
 * Date: 2025-12-11
 */

module config_regs (
    input  wire        clk,
    input  wire        rst_n,
    
    // Register Interface
    input  wire        reg_write,
    input  wire [3:0]  reg_addr, // 4-bit address for few registers
    input  wire [31:0] reg_wdata,
    output wire [31:0] reg_rdata,
    
    // Hardware Interface (To Controller)
    output reg         start,
    input  wire        done,
    
    output reg  [3:0]  kernel_h,
    output reg  [3:0]  kernel_w,
    output reg  [7:0]  input_h,
    output reg  [7:0]  input_w,
    output reg  [3:0]  stride,
    output reg  [3:0]  padding,
    output reg  [7:0]  output_h,
    output reg  [7:0]  output_w,
    output reg  [7:0]  input_channels,   // Total input channels
    output reg  [7:0]  output_channels  // Total output channels
);

    // Internal storage
    reg [31:0] ctrl_reg;
    // status_reg is purely combinational from inputs
    reg [31:0] kernel_dim_reg;
    reg [31:0] input_dim_reg;
    reg [31:0] param_reg;
    reg [31:0] output_dim_reg;
    reg [31:0] channel_reg;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            ctrl_reg       <= 0;
            kernel_dim_reg <= 0;
            input_dim_reg  <= 0;
            param_reg      <= 0;
            output_dim_reg <= 0;
            channel_reg    <= 0;
            
            start    <= 0;
            kernel_h <= 0;
            kernel_w <= 0;
            input_h  <= 0;
            input_w  <= 0;
            stride   <= 0;
            padding  <= 0;
            output_h <= 0;
            output_w <= 0;
            input_channels <= 16;   // Default 16
            output_channels <= 16;  // Default 16
        end else begin
            // Auto-clear start after 1 cycle (Pulse)
            if (start) start <= 0;
            
            if (reg_write) begin
                case (reg_addr)
                    4'h0: begin // Control
                        if (reg_wdata[0]) start <= 1;
                    end
                    // 4'h1: Status is RO
                    4'h2: begin // Kernel Dims (Addr 0x08 -> Index 2 if word addressed, let's assume byte addr >> 2)
                        kernel_dim_reg <= reg_wdata;
                        kernel_w <= reg_wdata[3:0];
                        kernel_h <= reg_wdata[11:8];
                    end
                    4'h3: begin // Input Dims (Addr 0x0C -> Index 3)
                        input_dim_reg <= reg_wdata;
                        input_w <= reg_wdata[7:0];
                        input_h <= reg_wdata[15:8];
                    end
                    4'h4: begin // Stride & Padding (Addr 0x10 -> Index 4)
                        param_reg <= reg_wdata;
                        stride    <= reg_wdata[3:0];
                        padding   <= reg_wdata[7:4];
                    end
                    4'h5: begin // Output Dims (Addr 0x14 -> Index 5)
                        output_dim_reg <= reg_wdata;
                        output_w <= reg_wdata[7:0];
                        output_h <= reg_wdata[15:8];
                    end
                    4'h6: begin // Channel Config (Addr 0x18 -> Index 6)
                        channel_reg <= reg_wdata;
                        input_channels <= reg_wdata[7:0];
                        output_channels <= reg_wdata[15:8];
                    end
                endcase
            end
        end
    end
    
    // Read Logic
    reg [31:0] reg_rdata_comb;
    always @(*) begin
        case (reg_addr)
            4'h0: reg_rdata_comb = {31'b0, start}; // Reflects current state
            4'h1: reg_rdata_comb = {31'b0, done};
            4'h2: reg_rdata_comb = kernel_dim_reg;
            4'h3: reg_rdata_comb = input_dim_reg;
            4'h4: reg_rdata_comb = param_reg;
            4'h5: reg_rdata_comb = output_dim_reg;
            4'h6: reg_rdata_comb = channel_reg;
            default: reg_rdata_comb = 32'd0;
        endcase
    end
    
    assign reg_rdata = reg_rdata_comb;

endmodule
